      --
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package tipos is

type ESTADOS is (F, ID, EX, MEM, WB);

type matrix is array(0 to 15) of std_logic_vector(0 to 7);

constant DOSPUNTOS: matrix:=(
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00011100",
"00011100",
"00011100",
"00000000",
"00000000",
"00000000",
"00011100",
"00011100",
"00011100",
"00000000"
);

constant VACIO: matrix:=(
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000"
);
constant CERO: matrix:=(
"00000000",
"01111110",
"01111110",
"01111110",
"01000010",
"01000010",
"01000010",
"01000010",
"01000010",
"01000010",
"01000010",
"01000010",
"01111110",
"01111110",
"01111110",
"00000000"
);
constant UNO: matrix:=(
"00000000",
"01111110",
"01111110",
"01111110",
"01111110",
"01111110",
"01111110",
"01111110",
"01111110",
"01111110",
"01111110",
"01111110",
"01111110",
"01111110",
"01111110",
"00000000"
);

constant A: matrix:=(
"00000000",
"00111100",
"00111100",
"01111110",
"01100110",
"01100110",
"01100110",
"01100110",
"01111110",
"01111110",
"01111110",
"01100110",
"01100110",
"01100110",
"01100110",
"00000000"
);

constant B: matrix:=(
"00000000",
"01111100",
"01111110",
"01100110",
"01100110",
"01100110",
"01100100",
"01111100",
"01111100",
"01100100",
"01100110",
"01100110",
"01100110",
"01111110",
"01111100",
"00000000"
);

constant C: matrix:=(
"00000000",
"00111110",
"01111110",
"01100000",
"01100000",
"01100000",
"01100000",
"01100000",
"01100000",
"01100000",
"01100000",
"01100000",
"01100000",
"01111110",
"00111110",
"00000000"
);

constant E: matrix:=(
"00000000",
"01111110",
"01111110",
"01100000",
"01100000",
"01100000",
"01100000",
"01111110",
"01111110",
"01100000",
"01100000",
"01100000",
"01100000",
"01111110",
"01111110",
"00000000"
);

constant FF: matrix:=(
"00000000",
"01111110",
"01111110",
"01100000",
"01100000",
"01100000",
"01100000",
"01111100",
"01111100",
"01100000",
"01100000",
"01100000",
"01100000",
"01100000",
"01100000",
"00000000"
);

constant D: matrix:=(
"00000000",
"01110000",
"01111000",
"01101100",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01101100",
"01111000",
"01110000",
"00000000"
);

constant G: matrix:=(
"00000000",
"00111110",
"01111110",
"01100000",
"01100000",
"01100000",
"01100000",
"01100000",
"01101110",
"01101110",
"01100110",
"01100110",
"01100110",
"01111110",
"00111100",
"00000000"
);

constant I: matrix:=(
"00000000",
"00011000",
"00011000",
"00000000",
"00000000",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00000000"
);

constant II: matrix:=(
"00000000",
"01111110",
"01111110",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"01111110",
"01111110",
"00000000"
);

constant J: matrix:=(
"00000000",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"01100110",
"01100110",
"01100110",
"01111110",
"00111100",
"00000000"
);

constant L: matrix:=(
"00000000",
"01100000",
"01100000",
"01100000",
"01100000",
"01100000",
"01100000",
"01100000",
"01100000",
"01100000",
"01100110",
"01100110",
"01100110",
"01111110",
"01111110",
"00000000"
);

constant N: matrix:=(
"00000000",
"01000010",
"01100010",
"01100010",
"01100010",
"01010010",
"01010010",
"01010010",
"01001010",
"01001010",
"01001010",
"01000110",
"01000110",
"01000110",
"01000010",
"00000000"
);

constant M: matrix:=(
"00000000",
"01000010",
"01100110",
"01100110",
"01100110",
"01011010",
"01011010",
"01011010",
"01000010",
"01000010",
"01000010",
"01000010",
"01000010",
"01000010",
"01000010",
"00000000"
);

--constant NN: matrix:=(
--"00000000",
--"00011000",
--"00100100",
--"01000010",
--"01000010",
--"01000010",
--"01000010",
--"01000010",
--"01000010",
--"01000010",
--"01000010",
--"01000010",
--"01000010",
--"01000010",
--"01000010",
--"00000000"
--);


constant O: matrix:=(
"00000000",
"00111100",
"01111110",
"01111110",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01111110",
"01111110",
"00111100",
"00000000"
);

constant P: matrix:=(
"00000000",
"00111100",
"01111110",
"01100110",
"01100110",
"01100110",
"01100110",
"01111110",
"01111100",
"01100000",
"01100000",
"01100000",
"01100000",
"01100000",
"01100000",
"00000000"
);

constant Q: matrix:=(
"00000000",
"00111100",
"01111110",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01111110",
"00111100",
"00001100",
"00000110",
"00000000"
);

constant R: matrix:=(--no me gusta
"00000000",
"00111100",
"01111110",
"01100110",
"01100110",
"01100110",
"01100100",
"01111100",
"01111100",
"01100100",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"00000000"
);

constant S: matrix:=(
"00000000",
"00111110",
"01111110",
"01100000",
"01100000",
"01100000",
"01100000",
"01111100",
"01111110",
"00000110",
"00000110",
"00000110",
"00000110",
"01111110",
"01111100",
"00000000"
);

constant T: matrix:=(
"00000000",
"01111110",
"01111110",
"01111110",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00011000",
"00000000"
);

constant U: matrix:=(
"00000000",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01100110",
"01111110",
"01111110",
"00111100",
"00000000"
);

constant W: matrix:=(
"00000000",
"01000100",
"01000100",
"01000100",
"01000100",
"01000100",
"01000100",
"01000100",
"01000100",
"01010100",
"01010100",
"01010100",
"01111100",
"01111100",
"01101100",
"00000000"
);

constant X: matrix:=(
"00000000",
"01000010",
"01000010",
"01000010",
"00100100",
"00100100",
"00100100",
"00011000",
"00011000",
"00100100",
"00100100",
"00100100",
"01000010",
"01000010",
"01000010",
"00000000"
);

end tipos;

package body tipos is


 
end tipos;